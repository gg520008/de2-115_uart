library verilog;
use verilog.vl_types.all;
entity diven_vlg_check_tst is
    port(
        diven           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end diven_vlg_check_tst;
