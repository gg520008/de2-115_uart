library verilog;
use verilog.vl_types.all;
entity fifo_vlg_vec_tst is
end fifo_vlg_vec_tst;
