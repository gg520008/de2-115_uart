library verilog;
use verilog.vl_types.all;
entity diven_vlg_vec_tst is
end diven_vlg_vec_tst;
