library verilog;
use verilog.vl_types.all;
entity mydelay_vlg_vec_tst is
end mydelay_vlg_vec_tst;
