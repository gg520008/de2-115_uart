library verilog;
use verilog.vl_types.all;
entity uart_top_tf is
end uart_top_tf;
